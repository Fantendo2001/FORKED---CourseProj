`timescale 1ns/1ps

module alu_test;

reg[31:0] a,b;
reg[15:0] immediate;
reg[4:0] opcode;

wire[31:0] c, HI, LO;
wire zero;
wire overflow;
wire neg;

parameter  sla = 5'b00000,
srai = 5'b00001,
add = 5'b00010,
sub = 5'b00011,
mult = 5'b00100,
div = 5'b00101,
addi = 5'b00110,
addu = 5'b00111,
subu = 5'b01000,
multu = 5'b01001,
divu = 5'b01010,
addiu = 5'b01011,
sqrt = 5'b01100,
_and = 5'b01101,
_or = 5'b01110,
_nor = 5'b01111,
_xor = 5'b10000,
_xnor = 5'b10001,
andi = 5'b10010,
ori = 5'b10011,
slt = 5'b10100,
slti = 5'b10101;

alu testalu(a,b,immediate,opcode,c,HI,LO,zero,overflow,neg);


initial
begin

$display("op: a      : b      : imm: c      : HI     : LO     : zf: of: nf: reg_A  : reg_B  : reg_C");
$monitor(" %h:%h:%h:%h:%h:%h:%h: %h : %h : %h :%h:%h:%h",
opcode, a, b, immediate, c, HI, LO, zero, overflow, neg, testalu.reg_A, testalu.reg_B, testalu.reg_C);

//// arith left shift

#10 a=32'b1101_1101_1101_1101_1101_1101_1101_1101;
opcode= sla;//5'b00000

#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
opcode= sla;


//// arith right shift

#10 a=32'b1111_1101_1111_1101_1111_1101_1111_1101;
opcode= srai; //5'b00001

#10 a=32'b0011_1001_0011_1001_0011_1001_0011_1001;
opcode= srai;

//// add

#10 a=32'b1000_0000_0000_0000_0000_0000_0000_0000;
    b=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    opcode = add;

//// sub

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    b=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    opcode = sub;

//// mult

#10 a=32'b1000_0000_0000_0000_0000_0000_0000_0010;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    opcode = mult;

//// div

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    opcode = div;

//// addi

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    immediate=16'b1111_1111_1111_1111;
    opcode = addi;

//// addu

#10 a=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    b=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    opcode = addu;

//// subu

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    b=32'b1000_0000_0000_0000_0000_0000_0000_0000;
    opcode = subu;


//// multu

#10 a=32'b1000_0000_0000_0000_0000_0000_0000_0010;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    opcode = multu;


//// divu

#10 a=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    b=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    opcode = divu;


//// addiu

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    immediate=16'b1111_1111_1111_1111;
    opcode = addiu;


//// _and

#10 a=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    b=32'b1111_1111_0000_1111_0000_1111_0000_1111;
    opcode = _and;


//// _or

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    opcode = _or;


//// _nor

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    opcode = _nor;


//// _xor

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    opcode = _xor;


//// _xnor

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    opcode = _xnor;


//// andi

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    immediate=16'b1111_1111_1111_1111;
    opcode = andi;


//// ori

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    immediate=16'b1111_1111_1111_1111;
    opcode = ori;


//// slt

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    opcode = slt;


//// slti

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    b=16'b0000_0000_0000_0111;
    opcode = slti;


#10 $finish;
end
endmodule


